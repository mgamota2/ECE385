module LEDvect(	input [15:0] IR,
						input LD_LED, Clk,
						output [9:0] LED

);

	
	
endmodule