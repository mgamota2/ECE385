module mp_toplevel(
	input logic Clk, Run, Continue,
	input logic [9:0] SW,
	output logic [9:0] LED,
	output logic [6:0] HEX0, HEX1, HEX2, HEX3

);

endmodule