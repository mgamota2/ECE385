//------------------------------------------------------------------------------
// Company:          UIUC ECE Dept.
// Engineer:         Stephen Kempf
//
// Create Date:    17:44:03 10/08/06
// Design Name:    ECE 385 Lab 6 Given Code - Incomplete ISDU
// Module Name:    ISDU - Behavioral
//
// Comments:
//    Revised 03-22-2007
//    Spring 2007 Distribution
//    Revised 07-26-2013
//    Spring 2015 Distribution
//    Revised 02-13-2017
//    Spring 2017 Distribution
//------------------------------------------------------------------------------
`include "SLC3_2.sv"
import SLC3_2::*;

module ISDU (   input logic         Clk, 
									Reset,
									Run,
									Continue,
									
				input logic[3:0]    Opcode, 
				input logic         IR_5,
				input logic         IR_11,
				input logic         BEN,
				  
				output logic        LD_MAR,
									LD_MDR,
									LD_IR,
									LD_BEN,
									LD_CC,
									LD_REG,
									LD_PC,
									LD_LED, // for PAUSE instruction
									
				output logic        GatePC,
									GateMDR,
									GateALU,
									GateMARMUX,
									
				output logic [1:0]  PCMUX,
				output logic        DRMUX,
									SR1MUX,
									SR2MUX,
									ADDR1MUX,
				output logic [1:0]  ADDR2MUX,
									ALUK,
				  
				output logic        Mem_OE,
									Mem_WE
				);

//	enum logic [3:0] {  Halted, 
//						PauseIR1, 
//						PauseIR2, 
//						S_18, 
//						S_33_1, 
//						S_33_2,
//						S_33_3,
//						S_35, 
//						S_32, 
//						S_01}   State, Next_state;   // Internal state logic
						
	////Week 2
	enum logic [4:0] {S_01,S_5,S_9,S_6,S_25, S_25_1, S_25_2,S_27,S_7,S_23,S_16, S_16_1, S_16_2,
							S_21,S_4,S_12,S_22,S_18,S_33_1,S_33_2, S_33_3,
 						  S_35,S_32,S_0, PauseIR1, PauseIR2, Halted} State, Next_state;
		
	always_ff @ (posedge Clk)
	begin
		if (Reset) 
			State <= Halted;
		else 
			State <= Next_state;
	end
   
	always_comb
	begin 
		// Default next state is staying at current state
		Next_state = State;
		
		// Default controls signal values
		LD_MAR = 1'b0;
		LD_MDR = 1'b0;
		LD_IR = 1'b0;
		LD_BEN = 1'b0;
		LD_CC = 1'b0;
		LD_REG = 1'b0;
		LD_PC = 1'b0;
		LD_LED = 1'b0;
		 
		GatePC = 1'b0;
		GateMDR = 1'b0;
		GateALU = 1'b0;
		GateMARMUX = 1'b0;
		 
		ALUK = 2'b00;
		 
		PCMUX = 2'b00;
		DRMUX = 1'b0;
		SR1MUX = 1'b0;
		SR2MUX = 1'b0;
		ADDR1MUX = 1'b0;
		ADDR2MUX = 2'b00;
		 
		Mem_OE = 1'b0;
		Mem_WE = 1'b0;
	
		// Assign next state
		unique case (State)
			Halted : 
				if (Run) 
					Next_state = S_18;                      
			S_18 : 
				Next_state = S_33_1;
			// Any states involving SRAM require more than one clock cycles.
			// The exact number will be discussed in lecture.
			S_33_1 : 
				Next_state = S_33_2;
			S_33_2 : 
				Next_state = S_33_3;
			S_33_3 : 
				Next_state = S_35;
			S_35 : 
				Next_state = S_32;
			// PauseIR1 and PauseIR2 are only for Week 1 such that TAs can see 
			// the values in IR.
			PauseIR1 : 
				if (~Continue) 
					Next_state = PauseIR1;
				else 
					Next_state = PauseIR2;
			PauseIR2 : 
				if (Continue) 
					Next_state = PauseIR2;
				else 
					Next_state = S_18;
			S_32 : 
				case (Opcode)
					op_ADD : 
						Next_state = S_01;
					op_AND : 
						Next_state = S_5;
					op_NOT : 
						Next_state = S_9;
					op_LDR : 
						Next_state = S_6;
					op_STR : 
						Next_state = S_7;
					op_JSR : 
						Next_state = S_4;
					op_JMP : 
						Next_state = S_12;
					op_BR : 
						Next_state = S_0;
					op_PSE : 
						Next_state = PauseIR1;
					NO_OP : 
						Next_state = State;

					default : 
						Next_state = S_18;
				endcase
			//ADD
			S_01 : 
				Next_state = S_18;				
			//AND
			S_5 : 
				Next_state = S_18;
			//NOT
			S_9 : 
				Next_state = S_18;
			//LDR
			S_6 : 
				Next_state = S_25;
			S_25 : 
				Next_state = S_25_1;
			S_25_1 : 
				Next_state = S_25_2;
			S_25_2 : 
				Next_state = S_27;
			S_27 : 
				Next_state = S_18;
			//STR
			S_7 : 
				Next_state = S_23;
			S_23 : 
				Next_state = S_16;
			S_16 : 
				Next_state = S_16_1;
			S_16_1 : 
				Next_state = S_16_2;
			S_16_2 : 
				Next_state = S_18;
			//JSR
			S_4 : 
				Next_state = S_21;
			S_21 : 
				Next_state = S_18;
			//JMP
			S_12 : 
				Next_state = S_18;
			//BR
			S_0 : 
				if (BEN)
					Next_state = S_22;
				else
					Next_state = S_18;
			S_22:
				Next_state = S_18;
				

			

			default : ;

		endcase
		
		// Assign control signals based on current state
		case (State)
			Halted: ;
			S_18 : 
				begin 
					GatePC = 1'b1;
					LD_MAR = 1'b1;
					PCMUX = 2'b00;
					LD_PC = 1'b1;
				end
			S_33_1 : 
				Mem_OE = 1'b1;
			S_33_2 : 
				begin 
					Mem_OE = 1'b1;
					LD_MDR = 1'b1;
				end
			S_33_3 : 
				begin 
					Mem_OE = 1'b1;
					LD_MDR = 1'b1;
				end
			S_35 : 
				begin 
					GateMDR = 1'b1;
					LD_IR = 1'b1;
				end
			PauseIR1: ;
			PauseIR2: ;
			S_32 : 
				LD_BEN = 1'b1;
			S_01 : 
				begin 
					SR2MUX = IR_5;
					SR1MUX = 1'b1;
					DRMUX=1'b1;
					ALUK = 2'b00;
					GateALU = 1'b1;
					LD_REG = 1'b1;
					LD_CC=1'b1;
				end
			S_5:
				begin 
					SR2MUX = IR_5;
					SR1MUX = 1'b1;
					DRMUX=1'b1;
					ALUK = 2'b10;
					GateALU = 1'b1;
					LD_REG = 1'b1;
					LD_CC=1'b1;
				end
			S_9:
				begin 
					SR2MUX = 1'b0;
					SR1MUX = 1'b1;
					ALUK = 2'b01;
					DRMUX=1'b1;
					GateALU = 1'b1;
					LD_REG = 1'b1;
					LD_CC=1'b1;
				end
			S_6:
				begin
					GateMARMUX=1'b1;
					ADDR2MUX=2'b01;
					ADDR1MUX=1'b1;
					SR1MUX=1'b0;
					LD_MAR=1'b1;
					
				end
			S_25:
				begin
					Mem_OE=1'b1;
					LD_MDR=1'b1;					
				end
			S_27:
				begin
					GateMDR=1'b1;
					DRMUX=1'b1;
					LD_REG=1'b1;
					LD_CC=1'b1;
				end
			S_7:
				begin
					GateMARMUX=1'b1;
					ADDR2MUX=2'b01;
					ADDR1MUX=1'b1;
					SR1MUX=1'b0;
					LD_MAR=1'b1;
					
				end
			S_23:
				begin
					SR1MUX=1'b0;
					ADDR1MUX=1'b1;
					ADDR2MUX=2'b00;
					GateMARMUX=1'b1;
					Mem_OE=1'b0;
					LD_MDR=1'b1;
				end
			S_16:
				begin
					GateMDR=1'b1;
					LD_MAR=1'b1;
				end
			S_4:
				begin
					LD_REG=1'b1;
					GatePC=1'b1;
					DRMUX=1'b0;	
				end
			S_21:
				begin
					ADDR1MUX=1'b0;
					ADDR2MUX=2'b11;
					PCMUX=2'b01;
					LD_PC=1'b1;
				end
			S_12:
				begin
					PCMUX=2'b01;
					ADDR2MUX=2'b00;
					LD_PC=1'b1;
					SR1MUX=1'b1;
					ADDR1MUX=1'b1;
				end
			S_22:
				begin
					LD_PC=1'b1;
					ADDR1MUX=1'b0;
					PCMUX=2'b01;
					ADDR2MUX=2'b10;
				end
			

			// You need to finish the rest of states.....

			default : ;
		endcase
	end 

	
endmodule
